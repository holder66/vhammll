// load_settings_test.v
module vhammll

fn test_read_multiple_opts() {
	dump(read_multiple_opts('/Users/henryolders/use_vhammll/vhammll/src/testdata/2_class.opts')!)
}
