// save_settings.v

module vhamml
