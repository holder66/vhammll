// rank
module vhammll

import maps

struct RankValue {
mut:
	attr_indx  int
	rank_value i64
	bin_no     int
}

const rank_help = '
Description:
  "rank" rank orders a dataset\'s attributes in terms of ability 
to distinguish between classes; it takes into account class prevalences.

Usage: `v run main.v rank <options> <path_to_dataset_file>`

Example: `v run .main.v rank -b 3,6 -x -wr datasets/iris.tab`

Options: 
  -b --bins, eg, "3,6" specifies the lower and upper limits for the number 
      of slices or bins for continuous attributes [Options.bins]
  -x --exclude, exclude missing values from rank value calculations [Parameters.exclude_flag]
  -g --graph, produce a plot showing rank values vs number of bins for   
      continuous attributes [DisplaySettings.graph_flag]
  -l --limit-output, followed by an integer which specifies how many
  		attributes should be included in the console listing [DisplaySettings.limit_output]
  -of --overfitting, console output and graph to include information
  		allowing for an assessment of overfitting likelihood [DisplaySettings.overfitting_flag]
  -exr --explore-rank, followed by eg "2,7", will repeat the ranking
  		exercise over the binning range from 2 through 7 [Options.explore_rank]
  -u --uniform, uses uniform binning over all attributes [Parameters.uniform_bins]
  -wr, weight contribution to ranking by considering class 
      prevalences [Parameters.weight_ranking_flag]

    '

// rank_attributes takes a Dataset and returns a list of all the
// dataset's usable attributes, ranked in order of each attribute's
// ability to separate the classes.
// ```
// Algorithm:
// for each attribute:
// 	create a matrix with attribute values for row headers, and
// 	class values for column headers;
// 	for each unique value `val` for that attribute:
// 		for each unique value `class` of the class attribute:
// 			for each instance:
// 				accumulate a count for those instances whose class value
// 				equals `class`;
// 				populate the matrix with these accumulated counts;
// 	for each `val`:
// 		get the absolute values of the differences between accumulated
// 		counts for each pair of `class` values`;
// 		add those absolute differences;
// 	total those added absolute differences to get the raw rank value
// for that attribute.
// To obtain rank values weighted by class prevalences, use the same algorithm
// except before taking the difference of each pair of accumulated counts,
// multiply each count of the pair by the class prevalence of the other class.
// (Note: rank_attributes always uses class prevalences as weights)
//
// Obtain a maximum rank value by calculating a rank value for the class
// attribute itself.
//
// To obtain normalized rank values:
// for each attribute:
// 	divide its raw rank value by the maximum rank value and multiply by 100.
//
// Sort the attributes by descending rank values.
// ```
//
// ```sh
// Options:
// `binning`: specifies the range for binning (slicing) continous attributes;
// `weight_ranking_flag`: appplies prevalences of each class in calculating rankings;
// `exclude_flag`: exclude missing values when calculating rank values;
// `explore_rank`: gives start and end values for maximum binning number to be
//     over an exploration of ranking for different binning values;
//
// Output options:
// `show_flag`: print the ranked list to the console;
// `graph_flag`: generate plots of rank values for each attribute on the
//     y axis, with number of bins on the x axis.
// `overfitting_flag`: generates metrics/plots to help determine, for continuous
//     attributes, whether overfitting is occurring.
// `outputfile_path`: saves the result as json.
// ```
pub fn rank_attributes(ds Dataset, opts Options) RankingResult {
	mut result := RankingResult{
		LoadOptions:     ds.LoadOptions
		DisplaySettings: opts.DisplaySettings
		path:            ds.path
		// binning:                    get_binning(opts.bins)
		exclude_flag:               opts.exclude_flag
		weight_ranking_flag:        opts.weight_ranking_flag
		array_of_ranked_attributes: []RankedAttribute{cap: ds.useful_discrete_attributes.len +
			ds.useful_continuous_attributes.len}
	}
	mut binning := Binning{}
	if ds.useful_continuous_attributes.len != 0 {
		if opts.binning.lower > 0 {
			binning = opts.binning
		} else {
			binning = get_binning(opts.bins)
		}
	}
	result.binning = binning
	mut rank_value_map := map[int]i64{}
	mut binning_map := map[int]int{}
	mut rank_value_array_map := map[int][]i64{}
	mut highest_rank_value := i64(0) // as generated by the class attribute, used for normalizing other values
	// for each attribute in the dataset
	for i, _ in ds.attribute_names {
		// base action on whether the attribute is the class attribute, continuous, discrete, or to be ignored
		match true {
			i == ds.class_index {
				// rank the class attribute and use it to normalize the other rank values
				highest_rank_value = rank_discrete_attribute(i, ds, opts)
			}
			i in ds.useful_continuous_attributes.keys() {
				r_v, bin_number, rank_value_array := rank_continuous_attribute(i, ds,
					binning, opts.exclude_flag, opts.weight_ranking_flag, opts.overfitting_flag)
				rank_value_map[i] = r_v
				binning_map[i] = bin_number
				rank_value_array_map[i] = rank_value_array
			}
			i in ds.useful_discrete_attributes.keys() {
				rank_value_map[i] = rank_discrete_attribute(i, ds, opts)
			}
			else {}
		}
	}
	mut rank_values_array := maps.to_array(rank_value_map, fn (k int, v i64) RankValue {
		return RankValue{
			attr_indx:  k
			rank_value: v
		}
	})
	for mut rank_value in rank_values_array {
		rank_value.bin_no = binning_map[rank_value.attr_indx]
	}
	// custom sort on descending rank value, then ascending bins, then index
	custom_sort_fn := fn (a &RankValue, b &RankValue) int {
		if a.rank_value > b.rank_value {
			return -1
		}
		if a.rank_value < b.rank_value {
			return 1
		}
		if a.rank_value == b.rank_value {
			if a.bin_no > b.bin_no {
				return 1
			}
			if a.bin_no < b.bin_no {
				return -1
			}
			if a.bin_no == b.bin_no {
				if a.attr_indx < b.attr_indx {
					return -1
				}
				return 1
			}
			return 0
		}
		return 0
	}
	rank_values_array.sort_with_compare(custom_sort_fn)
	// rank_values_array.sort(a.rank_value > b.rank_value)
	for attr in rank_values_array {
		result.array_of_ranked_attributes << RankedAttribute{
			attribute_index:  attr.attr_indx
			attribute_name:   ds.attribute_names[attr.attr_indx]
			attribute_type:   ds.attribute_types[attr.attr_indx]
			rank_value:       f32(100.0 * f64(attr.rank_value) / highest_rank_value)
			rank_value_array: rank_value_array_map[attr.attr_indx].map(f32(100.0 * f64(it) / highest_rank_value)).reverse()
			bins:             attr.bin_no
		}
	}
	if (opts.show_flag || opts.expanded_flag) && opts.command == 'rank' {
		show_rank_attributes(result)
	}
	if opts.graph_flag && opts.command == 'rank' {
		plot_rank(result)
	}
	if opts.outputfile_path != '' {
		save_json_file[RankingResult](result, opts.outputfile_path)
	}
	return result
}

// get_rank_value_for_strings
fn get_rank_value_for_strings(values []string, class_values []string, class_counts map[string]int, opts Options) i64 {
	// println('values: $values  class_values: $class_values  class_counts: $class_counts')
	mut rank_val := i64(0)
	mut count := 0
	mut row := []int{}
	for unique_val, _ in element_counts(values) {
		if unique_val in opts.missings && opts.exclude_flag {
			continue
		}
		row = []int{}
		// loop through classes
		for class, _ in class_counts {
			// at this point, we have the columns and rows we need
			// now to populate it
			count = 0
			for i, val in values {
				if val == unique_val && class_values[i] == class {
					count += 1
				}
			}
			row << count
		}
		if opts.weight_ranking_flag {
			rank_val += sum_along_row_weighted(row, class_counts.values())
		} else {
			rank_val += sum_along_row_unweighted(row)
		}
	}
	return rank_val
}

// rank_discrete_attribute returns a rank value for attribute i.
fn rank_discrete_attribute(i int, ds Dataset, opts Options) int {
	mut weights := ds.class_counts.values()
	mut class_indices_by_case := []int{len: ds.class_values.len, init: find(ds.classes,
		ds.class_values[index])}
	case_values := if i == ds.class_index {
		ds.class_values
	} else {
		ds.useful_discrete_attributes[i]
	}
	uniques_values := uniques(case_values)
	mut hits := [][]int{len: ds.classes.len, init: []int{len: uniques_values.len}}
	for idx, case in case_values {
		if case in opts.missings && opts.exclude_flag {
			continue
		}
		uniques_index := find(uniques_values, case)
		hits[class_indices_by_case[idx]][uniques_index] += 1
	}
	return sum_absolute_differences(pairs(ds.classes.len), hits, weights, opts.weight_ranking_flag)
}

// rank_continuous_attribute calculates rank values for attribute i over a range of bin values given
// by opts.bins. It returns the maximum rank value found and the corresponding number of bins.
fn rank_continuous_attribute(i int, ds Dataset, binning_range Binning, exclude_flag bool, weight_ranking_flag bool, overfitting_flag bool) (int, int, []i64) {
	mut result := 0

	mut max_rank_value := 0
	mut bins_for_max_rank_value := 0
	mut rank_value_array := []i64{}
	values := ds.useful_continuous_attributes[i]
	mut weights := ds.class_counts.values()
	mut class_indices_by_case := []int{len: ds.class_values.len, init: find(ds.classes,
		ds.class_values[index])}
	for bin_number in binning_range.lower .. binning_range.upper + 1 {
		mut hits := [][]int{len: ds.classes.len, init: []int{len: bin_number + 1}}
		binning := discretize_attribute_with_range_check(values, array_min(values.filter(!is_nan(it))),
			array_max(values.filter(!is_nan(it))), bin_number)
		for j, val in binning {
			if val == 0 && exclude_flag {
				continue
			}
			hits[class_indices_by_case[j]][val] += 1
		}
		if overfitting_flag {
			dump('${i}    ${hits}')
		}
		// for each column in hits, sum up the absolute differences between each pair of values
		result = sum_absolute_differences(pairs(ds.classes.len), hits, weights, weight_ranking_flag)
		rank_value_array << result
		if result > max_rank_value {
			max_rank_value = result
			bins_for_max_rank_value = bin_number
		}
	}
	return max_rank_value, bins_for_max_rank_value, rank_value_array
}

// sum_absolute_differences sums up the absolute differences for each pair of entries in the hits list.
// if the weight_ranking_flag is set, the hits on either side of each pair are first multiplied by the
// prevalence of the class on the other side of the pair.
fn sum_absolute_differences(pair_values [][]int, hits [][]int, weights []int, weighting bool) int {
	mut rank_value := 0
	for k in pair_values {
		for m in 0 .. hits[0].len {
			if weighting {
				rank_value += abs_diff(hits[k[0]][m] * weights[k[1]], hits[k[1]][m] * weights[k[0]])
			} else {
				rank_value += abs_diff(hits[k[0]][m], hits[k[1]][m])
			}
		}
	}
	return rank_value
}

// sum_along_row_weighted returns the sum of the absolute values of
// the differences between counts multiplied by the class count for
// every combination pair of classes
fn sum_along_row_weighted(row []int, class_counts_array []int) i64 {
	mut row_sum := 0
	mut diff := 0
	for i, count1 in row#[..-1] {
		for j, count2 in row[i + 1..] {
			diff = count1 * class_counts_array[i + j + 1] - count2 * class_counts_array[i]
			// println('${i} ${j} ${count1} ${count2} ${class_counts_array[i + j + 1]} ${class_counts_array[i]}')
			if diff < 0 {
				diff *= -1
			}
			row_sum += diff
		}
	}
	// println('row_sum: $row_sum')
	return row_sum
}

// sum_along_row_unweighted returns the sum of the absolute values of
// the differences between counts
fn sum_along_row_unweighted(row []int) i64 {
	mut row_sum := 0
	mut diff := 0
	for i, count1 in row {
		for count2 in row[i + 1..] {
			diff = count1 - count2
			if diff < 0 {
				diff *= -1
			}
			row_sum += diff
		}
	}
	// println('row_sum: $row_sum')
	return row_sum
}

// abs_diff returns the absolute value of the difference between two numbers.
fn abs_diff[T](a T, b T) T {
	if a >= b {
		return a - b
	}
	return b - a
}

// pairs generates a list of permutations of the digits from 0 up to and including n, taken two at a time.
// Example: assert pairs(3) == [[0, 1], [0, 2], [1, 2]]
fn pairs(n int) [][]int {
	mut pair_list := [][]int{cap: n}
	for i in 0 .. n {
		for j in i + 1 .. n {
			pair_list << [i, j]
		}
	}
	return pair_list
}
