// main.v
module main
import vhamml

fn main() {
	vhamml.cli()!
}