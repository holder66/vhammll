module main

import vhammll

fn main() {
	vhammll.cli()!
}
