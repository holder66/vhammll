// save_settings.v

module vhammll
