// main.v
module main

import holder66.vhammll

fn main() {
	vhammll.cli()!
}
