// constants.v
module vhammll
