// show.v
// in order to establish style consistency, aim to use magenta underline
// for the first line of each output, and blue underline for table headings.
// use bold green for subheadings
// ie, println(m_u('\nfirst line')
// println(b_u('table header')
// println(g_b('subheading')
//
// this website https://towardsdatascience.com/multi-class-metrics-made-simple-part-ii-the-f1-score-ebe8b2c2ca1 gives the
// best explanation of multiclass metrics and how they're calculated

module vhammll

// import arrays
import strings
// import math

// pad
fn pad(l int) string {
	return strings.repeat(' '[0], l)
}

fn verbose_result(i int, cl Classifier, classify_result ClassifyResult) {
	println('case: ${i:-7}    classes: ${cl.classes.join(' | ')}')
	println('inferred class                   ratio    sphere index   radius   nearest neighbours')
	println('${classify_result.inferred_class:-30}  ${get_ratio(classify_result.nearest_neighbors_by_class):6.2f}    ${classify_result.sphere_index:12}   ${classify_result.hamming_distance:6}   ${classify_result.nearest_neighbors_by_class:-17}  \n')
}

// show_analyze prints out to the console, a series of tables detailing a
// dataset. It takes as input an AnalyzeResult struct generated by
// analyze_dataset().
pub fn show_analyze(result AnalyzeResult) {
	// println('result in show_analyze: ${result}')
	mut show := []string{}
	show << m_u('\nAnalysis of Dataset:') + lg(' ${result.datafile_path} ') +
		m('(File Type: ${result.datafile_type})')
	if result.class_missing_purge_flag {
		show << r('Note: instances with missing class values were purged.')
	}
	show << g_b('All Attributes:')
	show << b_u(' Index  Name${' ':36}Count  Uniques  Missing      %  Type')
	mut total_count := 0
	mut total_missings := 0

	for attr in result.attributes {
		show << '${attr.id:6}  ${attr.name:-37}  ${attr.count:6}  ${attr.uniques:7}  ${attr.missing:7}  ${attr.missing * 100 / f32(attr.count):5.1f}  ${attr.att_type:4}'
		total_count += attr.count
		total_missings += attr.missing
	}

	show << [
		'______${' ':40}_______           _______  _____',
		'Totals (less Class attribute)              ${total_count:10}        ${total_missings:10}  ${total_missings * 100 / f32(total_count):5.2f}%',
	]
	show << g_b('Counts of Attributes by Type')
	show << b_u('Type        Count')
	mut types := []string{}
	for attr in result.attributes {
		types << attr.att_type
	}
	for key, value in element_counts(types) {
		show << '${key}          ${value:6}'
	}
	show << 'Total:     ${types.len:6}'
	disc_atts := result.attributes.filter(it.for_training && it.att_type == 'D')
	show << g_b('Discrete Attributes for Training') + ' (${disc_atts.len} attributes)'
	show << b_u(' Index  Name${' ':34}Uniques  Missing      %')
	for attr in disc_atts {
		show << '${attr.id:6}  ${attr.name:-37} ${attr.uniques:7}  ${attr.missing:7}  ${attr.missing * 100 / f32(attr.count):5.1f}'
	}
	cont_atts := result.attributes.filter(it.for_training && it.att_type == 'C')
	show << g_b('Continuous Attributes for Training') + ' (${cont_atts.len} attributes)'

	show << b_u(' Index  Name${' ':34}Uniques  Missing      %        Min        Max' +
		'       Mean     Median')
	for attr in cont_atts {
		show <<
			'${attr.id:6}  ${attr.name:-37} ${attr.uniques:7}  ${attr.missing:7}  ${attr.missing * 100 / f32(attr.count):5.1f}' +
			' ${attr.min:10.3g} ${attr.max:10.3g} ${attr.mean:10.3g} ${attr.median:10.3g}'
	}
	show << g_b('The Class Attribute: "${result.class_name}"') +
		' (${result.class_counts.len} classes)'
	show << b_u('Class Value           Cases')
	for key, value in result.class_counts {
		show << '${key:-20}  ${value:5}'
	}
	print_array(show)
}

// show_rank_attributes prints to the console the ranked list of
// attributes in result, showing each attribute's name, index, type,
// rank value, and bin count. Output is limited to result.limit_output
// entries when that field is non-zero.
pub fn show_rank_attributes(result RankingResult) {
	mut exclude_phrase := 'included'
	if result.exclude_flag {
		exclude_phrase = 'excluded'
	}
	println(m_u('\nAttributes Sorted by Rank Value, for "${result.path}"'))
	println('Missing values: ${exclude_phrase}')
	println('Bin range for continuous attributes: from ${result.binning.lower} to ${result.binning.upper} with interval ${result.binning.interval}')
	println(if result.weight_ranking_flag { 'Weighted' } else { 'Unweighted' } +
		' by class prevalences')
	println('Purging of instances with missing class values: ${result.class_missing_purge_flag}')
	println(b_u('         Name                         Index  Type   Rank Value   Bins'))
	mut array_to_print := []string{}
	for i, attr in result.array_of_ranked_attributes {
		if result.limit_output != 0 && i >= result.limit_output {
			break
		}
		array_to_print << '${i + 1:6}   ${attr.attribute_name:-27} ${attr.attribute_index:6} ${attr.attribute_type:2}         ${attr.rank_value:7.2f} ${attr.bins:6}'
	}
	print_array(array_to_print)
}

// show_classifier outputs to the console information about a classifier
pub fn show_classifier(cl Classifier) {
	mut parameters_for_show := ParametersForShow{
		Parameters:  cl.Parameters
		LoadOptions: cl.LoadOptions
		Class:       cl.Class
	}
	println(m_u('\nClassifier from "${cl.datafile_path}"'))
	show_parameters(parameters_for_show)
	println(g_b('Trained attributes sorted by rank value:'))
	show_trained_attributes(cl.trained_attributes)
	println(g_b('\nClassifier History:'))
	println(b_u('Date & Time (UTC)    Event   From file                   Original Instances' +
		if cl.purge_flag { '  After purging' } else { '' }))
	// println(b_u('Date & Time (UTC)    Event   From file                   Original Instances  After purging',
	// 'underline'), 'blue'))
	for events in cl.history_events {
		println(
			'${events.event_date:-19}  ${events.event:-6}  ${events.file_path:-35} ${events.prepurge_instances_count:10}' +
			if cl.purge_flag { ' ${events.instances_count:14}' } else { '' })
	}
}

// show_parameters
fn show_parameters(r ParametersForShow) {
	if r.number_of_attributes.len == 1 {
		println('${'Number of attributes: ':55}' +
			if r.number_of_attributes[0] == 0 { 'all' } else { '${r.number_of_attributes[0]}' })
	}
	println('${'Binning range for continuous attributes: ':55}' +
		if r.binning.lower == 0 { 'not applicable (no continuous attributes used)' } else { 'from ${r.binning.lower} to ${r.binning.upper} with interval ${r.binning.interval}' })
	println('${'Missing values: ':55}' + if r.exclude_flag { 'excluded' } else { 'included' })
	println('${'Purging of duplicate instances: ':55}${r.purge_flag}')
	println('${'Prevalence weighting for ranking attributes: ':55}${r.weight_ranking_flag}')
	println('${'Prevalence weighting for nearest neighbor counts: ':55}${r.weighting_flag}')
	println('${'Add instances to balance class prevalences: ':55}${r.balance_prevalences_flag}')
	if r.balance_prevalences_flag {
		println('${'Threshold: ':60}${r.balance_prevalences_threshold}')
		println('${'class counts: ':60}${r.class_counts}   ratio: ${ratio(r.class_counts.values())}')
		println('${'pre_balance_prevalences_class_counts: ':60}${r.pre_balance_prevalences_class_counts}   ratio: ${ratio(r.pre_balance_prevalences_class_counts.values())}')
		// println('${'train_dataset_class_counts: ':60}${r.train_dataset_class_counts}   ratio: ${ratio(r.train_dataset_class_counts.values())}')
	}
	println('${'Purging of instances with missing class values: ':55}${r.class_missing_purge_flag}')
}

fn show_balanced_prevalences(load_options LoadOptions) {}

// show_validate prints to the console the results of a validate()
// run: the classifier parameters, the number of instances validated,
// and for each instance its index, inferred class, and nearest-
// neighbor counts by class.
pub fn show_validate(result ValidateResult) {
	mut parameters_for_show := ParametersForShow{
		Parameters:  result.Parameters
		LoadOptions: result.LoadOptions
		Class:       result.Class
	}
	println(m_u('\nValidation of "${result.validate_file_path}" using a classifier from "${result.datafile_path}"'))
	show_parameters(parameters_for_show)
	if result.purge_flag {
		total_count := result.prepurge_instances_counts_array[0]
		purged_count := total_count - result.classifier_instances_counts[0]
		purged_percent := 100 * f64(purged_count) / total_count
		println('Instances purged: ${purged_count} out of ${total_count} (${purged_percent:6.2f}%)')
	}
	println('Number of instances validated: ${result.inferred_classes.len}')
	println(c_u('  Index   Inferred Class    Nearest Neighbor Counts by Class (${result.classes})'))
	for i, val in result.inferred_classes {
		println('${i:7}   ${val:-14}    ${result.counts[i]}')
	}
}

// show_verify prints to the console the results of a verify() run:
// the classifier parameters (or multiple-classifier settings),
// instance counts, per-class accuracy, confusion matrix (when
// expanded), and binary metrics for two-class problems.
pub fn show_verify(result CrossVerifyResult, opts Options) {
	println(m_u('\nVerification of "${result.testfile_path}" using ' +
		if opts.multiple_flag { 'multiple classifiers ' } else { 'a classifier ' } +
		'from "${result.datafile_path}"'))
	if opts.multiple_flag {
		println('Classifier parameters are in file "${opts.multiple_classify_options_file_path}"')
		show_multiple_classifier_settings(result, opts)
	} else {
		mut parameters_for_show := ParametersForShow{
			Parameters:  result.Parameters
			LoadOptions: result.LoadOptions
			Class:       result.Class
		}
		show_parameters(parameters_for_show)
	}
	if result.purge_flag {
		total_count := result.prepurge_instances_counts_array[0]
		purged_count := total_count - result.classifier_instances_counts[0]
		purged_percent := 100 * f64(purged_count) / total_count
		println('Instances purged: ${purged_count} out of ${total_count} (${purged_percent:6.2f}%)')
	}
	if opts.show_attributes_flag {
		show_attributes_for_verify(result)
	}
	show_cross_or_verify_result(result, opts.DisplaySettings)
}

const headers = {
	0:  'Classifier ID:'
	1:  'Number of attributes:'
	2:  'Binning:'
	3:  'Exclude missing values:'
	4:  'Ranking using weighting:'
	5:  'Weighting of NN counts:'
	6:  'Balance prevalences:'
	7:  'Purge duplicate cases:'
	8:  'True / correct counts:'
	9:  'False / incorrect counts:'
	10: 'Raw accuracy:'
	11: 'Balanced accuracy:'
	12: 'Matthews Correlation Coef:'
	13: 'Sensitivity:'
	14: 'Specificity:'
	15: 'Maximum Hamming Distance:'
}

const attribute_headings = {
	0: '               Attribute:   '
	1: '  Index  RankValue  Bins:   '
}

// show_multiple_classifier_settings expects the multiple classifiers to be in opts, and
// the classifier indices in result
fn show_multiple_classifier_settings(result CrossVerifyResult, opts Options) {
	println('break_on_all_flag: ${opts.break_on_all_flag}     multi_strategy: ${opts.multi_strategy}     class_missing_purge_flag: ${opts.class_missing_purge_flag}')
	println(g_b('Multiple Classifier Parameters:'))
	show_multiple_classifier_settings_details(result.multiple_classifier_settings)
	if opts.show_attributes_flag {
		if result.multiple_classifier_settings.len > 0 {
			if opts.command == 'cross' {
				println(g_b('As trained attributes change from one fold to the next, they are not displayed for cross-validation operations.'))
			} else {
				// show_trained_attributes_for_multiple_classifier_settings(result.multiple_classifier_settings, result.classifier_indices)
			}
		} else {
			println(g_b('Unable to display Trained Attributes!'))
		}
	}
}

const minimum_column_width = 13

// show_multiple_classifier_settings_details displays on the console the parameters for each
// classifier used in a multiple classifier situation.
// the first parameter contains only the parameters for the classifiers to be displayed; the
// second parameter contains the classifier number to be shown.
// Returns an integer array with column widths.
fn show_multiple_classifier_settings_details(multiple_classifier_settings []ClassifierSettings) []int {
	if multiple_classifier_settings.len == 0 {
		println('Error Exit: multiple_classifier_settings in show_multiple_classifier_settings_details is empty')
		exit(1)
	}
	mut row_data := []string{len: headers.len, init: ''}
	mut col_width_array := []int{}
	for par in multiple_classifier_settings {
		a := par.Parameters
		b := par.BinaryMetrics
		c := par.Metrics
		d := par.LoadOptions
		corrects := c.correct_counts.map(it.str()).join(' ')
		incorrects := c.incorrect_counts.map(it.str()).join(' ')
		mut col_width := array_max([corrects.len, incorrects.len]) + 2
		if col_width < minimum_column_width {
			col_width = minimum_column_width
		}
		col_width_array << col_width
		row_data[0] += '${par.classifier_id:-13}' + pad(col_width - 13)
		row_data[1] += '${a.number_of_attributes[0]:-13}' + pad(col_width - 13)
		binning := '${a.binning.lower}, ${a.binning.upper}, ${a.binning.interval}'
		row_data[2] += '${binning:-13}' + pad(col_width - 13)
		row_data[3] += '${a.exclude_flag:-13}' + pad(col_width - 13)
		row_data[4] += '${a.weight_ranking_flag:-13}' + pad(col_width - 13)
		row_data[5] += '${a.weighting_flag:-13}' + pad(col_width - 13)
		row_data[6] += '${d.balance_prevalences_flag:-13}' + pad(col_width - 13)
		row_data[7] += '${a.purge_flag:-13}' + pad(col_width - 13)
		if c.class_counts_int.len > 2 {
			row_data[8] += corrects + pad(col_width - corrects.len)
			row_data[9] += incorrects + pad(col_width - incorrects.len)
			row_data[10] += '${b.raw_acc:-6.2f}%      ' + pad(col_width - 13)
			row_data[11] += '${c.balanced_accuracy:-6.2f}%      ' + pad(col_width - 13)
		} else {
			row_data[8] += '${b.t_p:-6} ${b.t_n:-6}' + pad(col_width - 13)
			row_data[9] += '${b.f_n:-6} ${b.f_p:-6}' + pad(col_width - 13)
			row_data[10] += '${b.raw_acc:-6.2f}%      ' + pad(col_width - 13)
			row_data[11] += '${b.bal_acc:-6.2f}%      ' + pad(col_width - 13)
			row_data[12] += '${b.mcc:-4.3f}        ' + pad(col_width - 13)
			row_data[13] += '${b.sens:-4.3f}        ' + pad(col_width - 13)
			row_data[14] += '${b.spec:-4.3f}        ' + pad(col_width - 13)
		}
		row_data[15] += '${a.maximum_hamming_distance:-13}' + pad(col_width - 13)
	}
	for i, row in row_data {
		if row != '' {
			println('${headers[i]:26}   ${row}')
		}
	}
	return col_width_array
}

// show_crossvalidation prints to the console the results of a
// cross_validate() run: the partitioning scheme, classifier
// parameters (or multiple-classifier settings), instance counts,
// per-class accuracy, confusion matrix (when expanded), and binary
// metrics for two-class problems.
pub fn show_crossvalidation(result CrossVerifyResult, opts Options) {
	println(m_u('\nCross-validation of "${result.datafile_path}"' +
		if opts.multiple_flag { ' using multiple classifiers' } else { '' }))
	println('Partitioning: ' + if result.folds == 0 { 'leave-one-out' } else { '${result.folds}-fold' + if result.repetitions > 1 { ', ${result.repetitions} repetitions' + if result.random_pick { ' with random selection of instances' } else { '' }
		 } else { ''
		 }
	 })
	if opts.multiple_flag {
		println('Classifier parameters are in file "${opts.multiple_classify_options_file_path}"')
		show_multiple_classifier_settings(result, opts)
	} else {
		mut parameters_for_show := ParametersForShow{
			Parameters:  result.Parameters
			LoadOptions: result.LoadOptions
			Class:       result.Class
		}
		show_parameters(parameters_for_show)
	}
	// if result.purge_flag {
	// 	total_count_avg := array_sum(result.prepurge_instances_counts_array) / f64(result.prepurge_instances_counts_array.len)
	// 	purged_count_avg := total_count_avg - array_sum(result.classifier_instances_counts) / f64(result.classifier_instances_counts.len)
	// 	purged_percent := 100 * purged_count_avg / total_count_avg
	// 	println('Average instances purged: ${purged_count_avg:10.1f} out of ${total_count_avg} (${purged_percent:6.2f}%)')
	// }
	// if opts.show_attributes_flag && !opts.multiple_flag && result.trained_attribute_maps_array.len > 0 {
	// 	println(g_b('Trained Attributes:'))
	// 	show_trained_attributes(result, [13])
	// } else {
	// 	println(g_b('Unable to display Trained Attributes!'))
	// }
	show_cross_or_verify_result(result, opts.DisplaySettings)
}

// show_cross_or_verify_result
fn show_cross_or_verify_result(result CrossVerifyResult, disp DisplaySettings) {
	println(g_b('Results:'))
	// mut metrics := get_metrics(result)
	if !disp.expanded_flag {
		percent := (f32(result.correct_count) * 100 / result.labeled_classes.len)
		println('correct inferences: ${result.correct_count} out of ${result.labeled_classes.len} (accuracy: raw:${percent:6.2f}% balanced:${result.balanced_accuracy:6.2f}%)')
	} else {
		show_expanded_result(result)
		print_confusion_matrix(result)
	}
}

// show_expanded_result
fn show_expanded_result(result CrossVerifyResult) {
	println(g('    Class                     Instances    True Positives    Precision    Recall    F1 Score'))
	show_multiple_classes_stats(result)
	if result.class_counts.len == 2 {
		println('A correct classification to "${result.pos_neg_classes[0]}" is a True Positive (TP);\nA correct classification to "${result.pos_neg_classes[1]}" is a True Negative (TN).')
		println("   TP    FN    TN    FP  Sens'y Spec'y    PPV    NPV  F1 Score  Accuracy: Raw  Balanced     MCC")
		println('${get_binary_stats_line(result)}')
	}
}

// get_show_bins
fn get_show_bins(bins []int) string {
	if bins == [] || 0 in bins {
		return '       '
	}
	if bins.len == 1 || bins[0] == bins[1] {
		return '${bins[0]:7}'
	}
	return '${bins[0]:2} - ${bins[1]:-2}'
}

// show_bins_for_trailer
fn show_bins_for_trailer(bins []int) string {
	if bins == [] || 0 in bins {
		return ''
	}
	if bins.len == 1 || bins[0] == bins[1] {
		return '${bins[0]}'
	}
	return '${bins[0]} - ${bins[1]}'
}

// print_confusion_matrix
fn print_confusion_matrix(result CrossVerifyResult) {
	// collect confusion matrix rows into a matrix
	mut confusion_matrix := [][]f64{}
	mut data_row := []f64{}
	for key, _ in result.confusion_matrix_map {
		data_row = []
		for _, value in result.confusion_matrix_map[key] {
			data_row << value
		}
		confusion_matrix << data_row
	}
	mut header_row := []string{}
	for key, _ in result.confusion_matrix_map {
		header_row << key
	}
	mut display_confusion_matrix := [][]string{}
	mut display_row := []string{}
	for row in confusion_matrix {
		display_row = []
		for col in row {
			display_row << '${col:10.1g}'
		}
		display_confusion_matrix << display_row
	}
	for i, class in header_row {
		display_confusion_matrix[i].prepend(class)
	}
	header_row.prepend('Predicted Classes (columns)')
	display_confusion_matrix.prepend([r('Actual Classes (rows)')])
	display_confusion_matrix.prepend(header_row)

	// get the length of the longest class name
	mut l := result.classes.map(it.len)
	l << 9 // to make sure that the minimum length covers up to 5 digits
	l_max := array_max(l)
	println(b_u('Confusion Matrix' +
		if result.repetitions > 1 { ' (values averaged over ${result.repetitions} repetitions):' } else { ':' }))
	mut padded_item := ''
	for i, rows in display_confusion_matrix {
		for j, item in rows {
			match true {
				i == 0 && j == 0 { // print first item in first row, ie 'predicted classes (columns)'
					print(r('${item}  '))
				}
				i == 0 { // print column headers, ie classes
					padded_item = '${pad(l_max - item.len + 2)}' + item
					print(c('${padded_item}'))
				}
				i == 1 && j == 0 { // print 'actual classes' header
					padded_item = '${pad(6)}' + item
					print(b('${padded_item}'))
				}
				j == 0 { // print first column (class names)
					padded_item = '${pad(27 - item.len)}' + item + '  '
					print(c('${padded_item}'))
				}
				else { // print numeric values for each cell
					padded_item = '${pad(l_max - item.len + 2)}' + item
					print('${padded_item}')
				}
			}
		}
		// carriage return at end of line
		println('')
	}
}

// get_binary_stats_line
fn get_binary_stats_line(r CrossVerifyResult) string {
	return '${r.t_p:5} ${r.f_n:5} ${r.t_n:5} ${r.f_p:5}   ${r.sens:5.3f}  ${r.spec:5.3f}  ${r.ppv:5.3f}  ${r.npv:5.3f}     ${r.f1_score_binary:5.3f}        ${r.raw_acc:6.2f}%   ${r.balanced_accuracy:6.2f}%   ${r.mcc:5.3f}'
}

// show_multiple_classes_stats
fn show_multiple_classes_stats(result CrossVerifyResult) {
	mut show_result := []string{}
	m := result.Metrics
	for i, class in result.classes {
		show_result << '    ${class:-27}   ${result.labeled_instances[class]:5}   ${result.correct_inferences[class]:5} (${f32(result.correct_inferences[class]) * 100 / result.labeled_instances[class]:6.2f}%)        ${m.precision[i]:5.3f}     ${m.recall[i]:5.3f}       ${m.f1_score[i]:5.3f}'
	}
	show_result << '        Totals                    ${result.total_count:5}   ${result.correct_count:5} (accuracy: raw:${result.raw_acc:6.2f}% balanced:${result.balanced_accuracy:6.2f}%)'
	for i, avg_type in m.avg_type {
		show_result << '${avg_type.title():20} Averages:                                   ${m.avg_precision[i]:5.3f}     ${m.avg_recall[i]:5.3f}       ${m.avg_f1_score[i]:5.3f}'
	}
	print_array(show_result)
}

// show_detailed_result
fn show_detailed_result(final_inferred_class string, labeled_classes []string, mcr MultipleClassifierResults) {
	println('classifier  sphere index  radius  nearest neighbors  ratio  inferred class')
	for i, icr in mcr.results_by_classifier {
		a := icr.results_by_radius.last()
		println('${mcr.classifiers[i]:10}  ${a.sphere_index:12}  ${a.radius:6}  ${a.nearest_neighbors_by_class:-17} ${get_ratio(a.nearest_neighbors_by_class):6.2f}  ${a.inferred_class} ')
	}
	println('           ${final_inferred_class} ${labeled_classes}')
}

// get_ratio
fn get_ratio(a []int) f64 {
	// println('a in get_ratio: ${a}')
	if a.all(it == 0) {
		return 1
	}
	if 0 in a {
		return f64(array_max(a.filter(it != 0)))
	}
	return f64(array_max(a)) / array_min(a)
}
