// save_settings.v

module hamml
